library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all; -- Package for arithmetic operations

----------------------------------------------------------
-- Entity declaration for clock enable
----------------------------------------------------------

entity clock_divider is
  generic (
    g_length : natural := 10 --! Length of a point in us. (500 000)
  );                       -- Note that there IS a semicolon between generic and port sections
  port (
    clk : in    std_logic; --! Main clock
    rst : in    std_logic; --! High-active synchronous reset
    ce  : out   std_logic  --! Clock enable pulse signal
  );
end entity clock_divider;

------------------------------------------------------------
-- Architecture body for clock enable
------------------------------------------------------------

architecture behavioral of clock_divider is

  -- Local counter
  signal sig_cnt : natural;

begin

  --------------------------------------------------------
  -- p_clk_enable:
  -- Generate clock enable signal. By default, enable signal
  -- is low and generated pulse is always one clock long.
  --------------------------------------------------------
  p_clk_divider : process (clk) is
  begin

    if rising_edge(clk) then                      -- Synchronous process
      if (rst = '1') then                         -- High-active reset
        sig_cnt <= 0;                             -- Clear local counter
        ce      <= '0';                           -- Set output to low

      -- Test number of clock periods
      elsif (sig_cnt = (g_length * 100 - 1)) then
        sig_cnt <= 0;                             -- Clear local counter
        ce      <= '1';                           -- Generate clock enable pulse
      else
        sig_cnt <= sig_cnt + 1;
        ce      <= '0';
      end if;
    end if;

  end process p_clk_divider;

end architecture behavioral;
